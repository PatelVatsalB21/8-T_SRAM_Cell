* c:\users\vatsal\8t_sram.cir
.lib "sky130_fd_pr/models/sky130.lib.spice" tt 


xm5 gnd writtenbit net-_m3-pad2_ gnd sky130_fd_pr__nfet_01v8
xm3 net-_m3-pad1_ net-_m3-pad2_ writtenbit net-_m3-pad1_ sky130_fd_pr__pfet_01v8
xm7 net-_m3-pad2_ writeenable bitbar gnd sky130_fd_pr__nfet_01v8
xm8 net-_m3-pad2_ bitbar net-_m8-pad3_ gnd sky130_fd_pr__nfet_01v8
xm4 gnd net-_m3-pad2_ writtenbit gnd sky130_fd_pr__nfet_01v8
xm1 writtenbit bitline net-_m1-pad3_ gnd sky130_fd_pr__nfet_01v8
xm2 writtenbit writeenable bitline gnd sky130_fd_pr__nfet_01v8
xm6 net-_m3-pad1_ writtenbit net-_m3-pad2_ net-_m3-pad1_ sky130_fd_pr__pfet_01v8
v5  net-_m8-pad3_ gnd 1.8
v2  writeenable gnd 1.8
v4  net-_m3-pad1_ gnd 1.8
v3  net-_m1-pad3_ gnd 1.8
* u1  writtenbit plot_v1
* u3  writeenable plot_v1
* u2  bitline plot_v1
* u4  bitbar plot_v1
v1  bitline gnd pulse(0v 1.8v 0u 0u 0u 10n 20n)
v6  bitbar gnd pulse(1.8v 0v 0u 0u 0u 10n 20n)
.tran 250e-12 20e-09 0e-06

* Control Statements 
.control
run
print allv > plot_data_v.txt
print alli > plot_data_i.txt
plot v(writtenbit)
plot v(writeenable)
plot v(bitline)
plot v(bitbar)
.endc
.end
